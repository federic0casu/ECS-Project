library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

package utilities is
        type arr is array(natural range <>) of std_logic_vector(7 downto 0);
end package;

package body utilities is 
end package body utilities;