library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

library work;
    use work.common_pkg.all;

entity full_adder_tree_tb is
end entity;

architecture architecture_of_tb of full_adder_tree_tb is
    -----------------------------------------------------------------------------------
    -- Testbench constants
    -----------------------------------------------------------------------------------
    constant T_CLK          : time     := 8 ns;   -- Clock period
    constant T_RESET        : time     := 100 ns; -- Period before the reset deassertion
    constant M_TB           : positive := 8;
    -----------------------------------------------------------------------------------
    -- End testbench constants
    -----------------------------------------------------------------------------------

    -----------------------------------------------------------------------------------
    -- Testbench signals
    -----------------------------------------------------------------------------------
    signal clk_tb       : std_logic := '0';  					
    signal arstn_tb     : std_logic := '0';  					
    signal enable_tb    : std_logic := '0';
    signal end_sim      : std_logic := '1';
    signal a_tb         : VECTOR(M_TB-1 downto 0);
    signal b_tb         : VECTOR(M_TB-1 downto 0);
    signal s_tb         : std_logic_vector(M_TB-1 downto 0);
    -----------------------------------------------------------------------------------
    -- End testbench signals
    -----------------------------------------------------------------------------------

    -----------------------------------------------------------------------------------
    -- Component to test (DUT) declaration
    -----------------------------------------------------------------------------------
    component full_adder_tree is
        generic (
            M    : positive
        );
        port (
            A   : in  VECTOR(M-1 downto 0);
            B   : in  VECTOR(M-1 downto 0);
            S   : out std_logic_vector(N_BIT-1 downto 0)
        );
    end component;
    -----------------------------------------------------------------------------------
    -- End component to test declaration
    -----------------------------------------------------------------------------------
begin

    DUT: full_adder_tree
        generic map (
            M => 8
        )
        port map (
            A => a_tb,
            B => b_tb,
            S => s_tb
        );

    clk_tb   <= not(clk_tb) and end_sim after T_CLK / 2; 
											                -- When end_sim is forced low, the clock stops toggling and the simulation ends.
    arstn_tb <= '1' after T_RESET;

    
    STIMULI : process(clk_tb, arstn_tb) 

        variable t : integer := 0;
        begin
            if (log2(M_TB) > 3 or log2(M_TB) < 3) then
                report "log2(M) = " & natural'image(log2(M_TB));
            elsif arstn_tb = '0' then
                t := 0;
                a_tb(0) <= "00000000"; 
                a_tb(1) <= "00000000"; 
                a_tb(2) <= "00000000"; 
                a_tb(3) <= "00000000";
                a_tb(4) <= "00000000"; 
                a_tb(5) <= "00000000"; 
                a_tb(6) <= "00000000"; 
                a_tb(7) <= "00000000";
            ------------------------------
                b_tb(0) <= "00000000"; 
                b_tb(1) <= "00000000"; 
                b_tb(2) <= "00000000"; 
                b_tb(3) <= "00000000";
                b_tb(4) <= "00000000"; 
                b_tb(5) <= "00000000"; 
                b_tb(6) <= "00000000"; 
                b_tb(7) <= "00000000";
            elsif rising_edge(clk_tb) then
                case(t) is  								-- Specifying the input_tb and end_sim depending on the value 
                    when 10000 => end_sim  <= '0';  		    -- This command stops the simulation when t = 10000
                    --------------------------------------------------------------------------------------------------------
                    -- Initial condition 
                    --------------------------------------------------------------------------------------------------------
                    when  1 => report "S must be '00000000' - S = " & std_logic'image(s_tb(7)) & std_logic'image(s_tb(6)) 
                                                                    & std_logic'image(s_tb(5)) & std_logic'image(s_tb(4))
                                                                    & std_logic'image(s_tb(3)) & std_logic'image(s_tb(2))
                                                                    & std_logic'image(s_tb(1)) & std_logic'image(s_tb(0));
                    --------------------------------------------------------------------------------------------------------
                    -- End initial condition 
                    --------------------------------------------------------------------------------------------------------

                    --------------------------------------------------------------------------------------------------------
                    -- 1st test
                    --------------------------------------------------------------------------------------------------------
                    when 1000 => a_tb(0) <= "00000010"; a_tb(1) <= "00000010"; a_tb(2) <= "00000010"; a_tb(3) <= "00000010";
                                 a_tb(4) <= "00000001"; a_tb(5) <= "00000001"; a_tb(6) <= "00000001"; a_tb(7) <= "00000001"; 
                               
                                 b_tb(0) <= "00000011"; b_tb(1) <= "00000011"; b_tb(2) <= "00000011"; b_tb(3) <= "00000011";
                                 b_tb(4) <= "00000010"; b_tb(5) <= "00000010"; b_tb(6) <= "00000010"; b_tb(7) <= "00000010";
                    when 1001 => report "S must be '00101000' - S = " & std_logic'image(s_tb(7)) & std_logic'image(s_tb(6)) 
                                                                      & std_logic'image(s_tb(5)) & std_logic'image(s_tb(4))
                                                                      & std_logic'image(s_tb(3)) & std_logic'image(s_tb(2))
                                                                      & std_logic'image(s_tb(1)) & std_logic'image(s_tb(0));
                    --------------------------------------------------------------------------------------------------------
                    -- End 1st test 
                    --------------------------------------------------------------------------------------------------------

                    --------------------------------------------------------------------------------------------------------
                    -- 2nd test 
                    --------------------------------------------------------------------------------------------------------
                    when 2000 => a_tb(0) <= "00000011"; a_tb(1) <= "00000010"; a_tb(2) <= "00000010"; a_tb(3) <= "00000010";
                                 a_tb(4) <= "00000010"; a_tb(5) <= "00000010"; a_tb(6) <= "00000010"; a_tb(7) <= "00000010"; 
                               
                                 b_tb(0) <= "00000010"; b_tb(1) <= "00000010"; b_tb(2) <= "00000010"; b_tb(3) <= "00000010";
                                 b_tb(4) <= "00000011"; b_tb(5) <= "00000010"; b_tb(6) <= "00000010"; b_tb(7) <= "00000010";
                    when 2001 => report "S must be '00100010' - S = " & std_logic'image(s_tb(7)) & std_logic'image(s_tb(6)) 
                                                                      & std_logic'image(s_tb(5)) & std_logic'image(s_tb(4))
                                                                      & std_logic'image(s_tb(3)) & std_logic'image(s_tb(2))
                                                                      & std_logic'image(s_tb(1)) & std_logic'image(s_tb(0)); 
                    --------------------------------------------------------------------------------------------------------
                    -- End 2nd test 
                    --------------------------------------------------------------------------------------------------------

                    --------------------------------------------------------------------------------------------------------
                    -- 3rd test
                    --------------------------------------------------------------------------------------------------------
                    when 3000 => a_tb(0) <= "00001010"; a_tb(1) <= "00001010"; a_tb(2) <= "00001010"; a_tb(3) <= "00001010";
                                 a_tb(4) <= "00001010"; a_tb(5) <= "00001010"; a_tb(6) <= "00001010"; a_tb(7) <= "00001010"; 
                               
                                 b_tb(0) <= "00010100"; b_tb(1) <= "00010100"; b_tb(2) <= "00010100"; b_tb(3) <= "00010100";
                                 b_tb(4) <= "00010100"; b_tb(5) <= "00010100"; b_tb(6) <= "00010100"; b_tb(7) <= "00010100";
                    when 3001 => report "S must be '11110000' - S = " & std_logic'image(s_tb(7)) & std_logic'image(s_tb(6)) 
                                                                      & std_logic'image(s_tb(5)) & std_logic'image(s_tb(4))
                                                                      & std_logic'image(s_tb(3)) & std_logic'image(s_tb(2))
                                                                      & std_logic'image(s_tb(1)) & std_logic'image(s_tb(0)); 
                    --------------------------------------------------------------------------------------------------------
                    -- End 3rd test 
                    --------------------------------------------------------------------------------------------------------

                    --------------------------------------------------------------------------------------------------------
                    -- 4th test
                    --------------------------------------------------------------------------------------------------------
                    when 4000 => a_tb(0) <= "00000001"; a_tb(1) <= "00000010"; a_tb(2) <= "00000011"; a_tb(3) <= "00000100";
                                 a_tb(4) <= "00000101"; a_tb(5) <= "00000110"; a_tb(6) <= "00000111"; a_tb(7) <= "00001000"; 
                               
                                 b_tb(0) <= "00000010"; b_tb(1) <= "00000101"; b_tb(2) <= "00000100"; b_tb(3) <= "00000011";
                                 b_tb(4) <= "00001010"; b_tb(5) <= "00001001"; b_tb(6) <= "00001000"; b_tb(7) <= "00010000";
                    when 4001 => report "S must be '01011101' - S = " & std_logic'image(s_tb(7)) & std_logic'image(s_tb(6)) 
                                                                      & std_logic'image(s_tb(5)) & std_logic'image(s_tb(4))
                                                                      & std_logic'image(s_tb(3)) & std_logic'image(s_tb(2))
                                                                      & std_logic'image(s_tb(1)) & std_logic'image(s_tb(0)); 
                    --------------------------------------------------------------------------------------------------------
                    -- End 4th test 
                    --------------------------------------------------------------------------------------------------------

                    --------------------------------------------------------------------------------------------------------
                    -- 5th test
                    --------------------------------------------------------------------------------------------------------
                    when 5000 => a_tb(0) <= "00100001"; a_tb(1) <= "00100010"; a_tb(2) <= "00100011"; a_tb(3) <= "01010101";
                                 a_tb(4) <= "00100101"; a_tb(5) <= "01100110"; a_tb(6) <= "00001111"; a_tb(7) <= "00101000"; 
                               
                                 b_tb(0) <= "10100010"; b_tb(1) <= "00010101"; b_tb(2) <= "00100100"; b_tb(3) <= "01001011";
                                 b_tb(4) <= "00001010"; b_tb(5) <= "01001001"; b_tb(6) <= "01001010"; b_tb(7) <= "00010100";
                    when 5001 => report "S must be '01010100' - S = " & std_logic'image(s_tb(7)) & std_logic'image(s_tb(6)) 
                                                                      & std_logic'image(s_tb(5)) & std_logic'image(s_tb(4))
                                                                      & std_logic'image(s_tb(3)) & std_logic'image(s_tb(2))
                                                                      & std_logic'image(s_tb(1)) & std_logic'image(s_tb(0)); 
                    --------------------------------------------------------------------------------------------------------
                    -- End 5th test 
                    --------------------------------------------------------------------------------------------------------
                    when others => null;                    -- Specifying that nothing happens in the other cases
                    end case;
                t := t + 1;  								             
            end if;
    end process;
end architecture;
